module vadd_ctrl(
  input clk, 
  input start
  output [9:0] addr
);


  always @(posedge clk) begin 
    if (start)
       
  end

endmodule
